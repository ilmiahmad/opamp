magic
tech sky130A
magscale 1 2
timestamp 1729224934
<< nmos >>
rect -189 -69 -29 131
rect 29 -69 189 131
<< ndiff >>
rect -247 119 -189 131
rect -247 -57 -235 119
rect -201 -57 -189 119
rect -247 -69 -189 -57
rect -29 119 29 131
rect -29 -57 -17 119
rect 17 -57 29 119
rect -29 -69 29 -57
rect 189 119 247 131
rect 189 -57 201 119
rect 235 -57 247 119
rect 189 -69 247 -57
<< ndiffc >>
rect -235 -57 -201 119
rect -17 -57 17 119
rect 201 -57 235 119
<< poly >>
rect -189 131 -29 157
rect 29 131 189 157
rect -189 -107 -29 -69
rect -189 -141 -173 -107
rect -45 -141 -29 -107
rect -189 -157 -29 -141
rect 29 -107 189 -69
rect 29 -141 45 -107
rect 173 -141 189 -107
rect 29 -157 189 -141
<< polycont >>
rect -173 -141 -45 -107
rect 45 -141 173 -107
<< locali >>
rect -235 119 -201 135
rect -235 -73 -201 -57
rect -17 119 17 135
rect -17 -73 17 -57
rect 201 119 235 135
rect 201 -73 235 -57
rect -189 -141 -173 -107
rect -45 -141 -29 -107
rect 29 -141 45 -107
rect 173 -141 189 -107
<< viali >>
rect -235 -57 -201 119
rect -17 -57 17 119
rect 201 -57 235 119
rect -173 -141 -45 -107
rect 45 -141 173 -107
<< metal1 >>
rect -241 119 -195 131
rect -241 -57 -235 119
rect -201 -57 -195 119
rect -241 -69 -195 -57
rect -23 119 23 131
rect -23 -57 -17 119
rect 17 -57 23 119
rect -23 -69 23 -57
rect 195 119 241 131
rect 195 -57 201 119
rect 235 -57 241 119
rect 195 -69 241 -57
rect -185 -107 -33 -101
rect -185 -141 -173 -107
rect -45 -141 -33 -107
rect -185 -147 -33 -141
rect 33 -107 185 -101
rect 33 -141 45 -107
rect 173 -141 185 -107
rect 33 -147 185 -141
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
