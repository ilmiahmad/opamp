magic
tech sky130A
magscale 1 2
timestamp 1729429965
<< nwell >>
rect -176 -1609 622 489
<< nsubdiff >>
rect -140 419 -80 453
rect 526 419 586 453
rect -140 393 -106 419
rect 552 393 586 419
rect -140 -1539 -106 -1517
rect 552 -1539 586 -1517
rect -140 -1573 -80 -1539
rect 526 -1573 586 -1539
<< nsubdiffcont >>
rect -80 419 526 453
rect -140 -1517 -106 393
rect 552 -1517 586 393
rect -80 -1573 526 -1539
<< poly >>
rect -56 381 36 397
rect -56 347 -40 381
rect -6 347 36 381
rect -56 332 36 347
rect 6 326 36 332
rect 410 381 502 397
rect 410 347 452 381
rect 486 347 502 381
rect 410 331 502 347
rect 410 325 440 331
rect -56 -119 36 -103
rect -56 -153 -40 -119
rect -6 -153 36 -119
rect -56 -168 36 -153
rect 6 -174 36 -168
rect 410 -119 502 -103
rect 410 -153 452 -119
rect 486 -153 502 -119
rect 410 -169 502 -153
rect 410 -174 440 -169
rect 94 -674 194 -426
rect 252 -674 352 -426
rect 6 -931 36 -926
rect -56 -947 36 -931
rect -56 -981 -40 -947
rect -6 -981 36 -947
rect -56 -996 36 -981
rect 410 -931 440 -926
rect 410 -947 502 -931
rect 410 -981 452 -947
rect 486 -981 502 -947
rect 410 -997 502 -981
rect 6 -1431 36 -1425
rect -56 -1447 36 -1431
rect -56 -1481 -40 -1447
rect -6 -1481 36 -1447
rect -56 -1496 36 -1481
rect 410 -1431 440 -1422
rect 410 -1447 502 -1431
rect 410 -1481 452 -1447
rect 486 -1481 502 -1447
rect 410 -1497 502 -1481
<< polycont >>
rect -40 347 -6 381
rect 452 347 486 381
rect -40 -153 -6 -119
rect 452 -153 486 -119
rect -40 -981 -6 -947
rect 452 -981 486 -947
rect -40 -1481 -6 -1447
rect 452 -1481 486 -1447
<< locali >>
rect -140 419 -80 453
rect 526 419 586 453
rect -140 393 -106 419
rect 552 393 586 419
rect -56 347 -40 381
rect -6 347 10 381
rect 436 347 452 381
rect 486 347 502 381
rect -40 303 -6 347
rect 452 304 486 347
rect -56 -153 -40 -119
rect -6 -153 10 -119
rect 436 -153 452 -119
rect 486 -153 502 -119
rect -40 -198 -6 -153
rect 452 -196 486 -153
rect -40 -947 -6 -904
rect 452 -947 486 -904
rect -56 -981 -40 -947
rect -6 -981 10 -947
rect 436 -981 452 -947
rect 486 -981 502 -947
rect -40 -1447 -6 -1404
rect 452 -1447 486 -1404
rect -56 -1481 -40 -1447
rect -6 -1481 10 -1447
rect 436 -1481 452 -1447
rect 486 -1481 502 -1447
rect -140 -1539 -106 -1517
rect 552 -1539 586 -1517
rect -140 -1573 -80 -1539
rect 526 -1573 586 -1539
<< viali >>
rect -40 347 -6 381
rect 452 347 486 381
rect -40 -153 -6 -119
rect 452 -153 486 -119
rect -40 -981 -6 -947
rect 452 -981 486 -947
rect -40 -1481 -6 -1447
rect 452 -1481 486 -1447
<< metal1 >>
rect -52 381 6 387
rect -52 347 -40 381
rect -6 347 6 381
rect -52 341 6 347
rect 440 381 498 387
rect 440 347 452 381
rect 486 347 498 381
rect 440 341 498 347
rect -46 300 6 341
rect 446 300 492 341
rect -46 288 91 300
rect -46 112 39 288
rect 91 112 101 288
rect 200 276 246 289
rect 355 288 492 300
rect -46 100 91 112
rect 187 100 197 276
rect 249 100 259 276
rect 345 112 355 288
rect 407 112 492 288
rect 355 100 492 112
rect 118 -24 170 62
rect 266 10 276 62
rect 328 10 338 62
rect 118 -76 328 -24
rect -52 -119 6 -113
rect -52 -153 -40 -119
rect -6 -153 6 -119
rect -52 -159 6 -153
rect -46 -200 6 -159
rect 108 -162 118 -110
rect 170 -162 180 -110
rect 276 -162 328 -76
rect 440 -119 498 -113
rect 440 -153 452 -119
rect 486 -153 498 -119
rect 440 -159 498 -153
rect 446 -200 493 -159
rect -46 -400 91 -200
rect 200 -212 246 -200
rect 187 -388 197 -212
rect 249 -388 259 -212
rect 200 -400 246 -388
rect 356 -400 493 -200
rect 42 -604 87 -400
rect 189 -491 195 -439
rect 247 -443 253 -439
rect 359 -443 404 -400
rect 247 -488 404 -443
rect 247 -491 253 -488
rect 191 -604 197 -600
rect 42 -649 197 -604
rect 42 -700 87 -649
rect 191 -652 197 -649
rect 249 -652 255 -600
rect 359 -700 404 -488
rect -46 -900 91 -700
rect 200 -712 246 -700
rect 187 -888 197 -712
rect 249 -888 259 -712
rect 356 -900 493 -700
rect -46 -941 0 -900
rect -52 -947 6 -941
rect -52 -981 -40 -947
rect -6 -981 6 -947
rect -52 -987 6 -981
rect 118 -1024 170 -938
rect 266 -990 276 -938
rect 328 -990 338 -938
rect 446 -941 492 -900
rect 440 -947 498 -941
rect 440 -981 452 -947
rect 486 -981 498 -947
rect 440 -987 498 -981
rect 118 -1076 328 -1024
rect 108 -1162 118 -1110
rect 170 -1162 180 -1110
rect 276 -1162 328 -1076
rect -46 -1212 91 -1200
rect 200 -1212 246 -1200
rect 355 -1212 492 -1200
rect -46 -1388 39 -1212
rect 91 -1388 101 -1212
rect 187 -1388 197 -1212
rect 249 -1388 259 -1212
rect 345 -1388 355 -1212
rect 407 -1388 492 -1212
rect -46 -1400 91 -1388
rect 200 -1400 246 -1388
rect 355 -1400 492 -1388
rect -46 -1441 0 -1400
rect 446 -1441 492 -1400
rect -52 -1447 6 -1441
rect -52 -1481 -40 -1447
rect -6 -1481 6 -1447
rect -52 -1487 6 -1481
rect 440 -1447 498 -1441
rect 440 -1481 452 -1447
rect 486 -1481 498 -1447
rect 440 -1487 498 -1481
<< via1 >>
rect 39 112 91 288
rect 197 100 249 276
rect 355 112 407 288
rect 276 10 328 62
rect 118 -162 170 -110
rect 197 -388 249 -212
rect 195 -491 247 -439
rect 197 -652 249 -600
rect 197 -888 249 -712
rect 276 -990 328 -938
rect 118 -1162 170 -1110
rect 39 -1388 91 -1212
rect 197 -1388 249 -1212
rect 355 -1388 407 -1212
<< metal2 >>
rect 39 288 91 298
rect 355 288 407 298
rect 39 102 91 112
rect 195 276 251 286
rect 40 -442 90 102
rect 355 102 407 112
rect 195 90 251 100
rect 276 62 328 72
rect 276 -24 328 10
rect 118 -76 328 -24
rect 118 -110 170 -76
rect 118 -172 170 -162
rect 195 -212 251 -202
rect 195 -398 251 -388
rect 195 -439 247 -433
rect 40 -487 195 -442
rect 40 -1202 90 -487
rect 195 -497 247 -491
rect 197 -600 249 -594
rect 356 -603 406 102
rect 249 -648 406 -603
rect 197 -658 249 -652
rect 195 -712 251 -702
rect 195 -898 251 -888
rect 276 -938 328 -928
rect 276 -1024 328 -990
rect 118 -1076 328 -1024
rect 118 -1110 170 -1076
rect 118 -1172 170 -1162
rect 356 -1202 406 -648
rect 39 -1212 91 -1202
rect 39 -1398 91 -1388
rect 195 -1212 251 -1202
rect 195 -1388 197 -1376
rect 249 -1388 251 -1376
rect 195 -1398 251 -1388
rect 355 -1212 407 -1202
rect 355 -1398 407 -1388
<< via2 >>
rect 195 100 197 276
rect 197 100 249 276
rect 249 100 251 276
rect 195 -388 197 -212
rect 197 -388 249 -212
rect 249 -388 251 -212
rect 195 -888 197 -712
rect 197 -888 249 -712
rect 249 -888 251 -712
rect 195 -1376 197 -1212
rect 197 -1376 249 -1212
rect 249 -1376 251 -1212
<< metal3 >>
rect 185 276 261 398
rect 185 100 195 276
rect 251 100 261 276
rect 185 -212 261 100
rect 185 -388 195 -212
rect 251 -388 261 -212
rect 185 -712 261 -388
rect 185 -888 195 -712
rect 251 -888 261 -712
rect 185 -1212 261 -888
rect 185 -1376 195 -1212
rect 251 -1376 261 -1212
rect 185 -1500 261 -1376
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729203764
transform 1 0 21 0 1 -1300
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729203764
transform 1 0 425 0 1 -300
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729203764
transform 1 0 21 0 1 -300
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729203764
transform 1 0 21 0 1 -800
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729203764
transform 1 0 21 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729203764
transform 1 0 425 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729203764
transform 1 0 425 0 1 -1300
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729203764
transform 1 0 425 0 1 -800
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_0
timestamp 1729196901
transform 1 0 223 0 1 -1300
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_1
timestamp 1729196901
transform 1 0 223 0 1 200
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_C6L7Y6  sky130_fd_pr__pfet_01v8_C6L7Y6_0
timestamp 1729197876
transform 1 0 223 0 1 -836
box -223 -164 223 198
use sky130_fd_pr__pfet_01v8_XLJ7Y8  sky130_fd_pr__pfet_01v8_XLJ7Y8_0
timestamp 1729197876
transform 1 0 223 0 1 -264
box -223 -198 223 164
<< labels >>
flabel nsubdiffcont 226 436 226 438 0 FreeSans 160 0 0 0 vdd
port 0 nsew
flabel metal2 60 -54 60 -52 0 FreeSans 160 0 0 0 d6
port 1 nsew
flabel metal2 386 -56 386 -54 0 FreeSans 160 0 0 0 d7
port 2 nsew
flabel metal3 226 12 226 14 0 FreeSans 160 0 0 0 d5
port 3 nsew
flabel metal1 144 -8 144 -6 0 FreeSans 160 0 0 0 vin
port 4 nsew
flabel metal2 306 -12 306 -10 0 FreeSans 160 0 0 0 vip
port 5 nsew
<< end >>
