magic
tech sky130A
magscale 1 2
timestamp 1729197478
<< nwell >>
rect -223 -200 223 200
<< pmos >>
rect -129 -100 -29 100
rect 29 -100 129 100
<< pdiff >>
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
<< pdiffc >>
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
<< poly >>
rect -119 181 -39 197
rect -119 164 -103 181
rect -129 147 -103 164
rect -55 164 -39 181
rect 39 181 119 197
rect 39 164 55 181
rect -55 147 -29 164
rect -129 100 -29 147
rect 29 147 55 164
rect 103 164 119 181
rect 103 147 129 164
rect 29 100 129 147
rect -129 -147 -29 -100
rect -129 -164 -103 -147
rect -119 -181 -103 -164
rect -55 -164 -29 -147
rect 29 -147 129 -100
rect 29 -164 55 -147
rect -55 -181 -39 -164
rect -119 -197 -39 -181
rect 39 -181 55 -164
rect 103 -164 129 -147
rect 103 -181 119 -164
rect 39 -197 119 -181
<< polycont >>
rect -103 147 -55 181
rect 55 147 103 181
rect -103 -181 -55 -147
rect 55 -181 103 -147
<< locali >>
rect -119 147 -113 181
rect -45 147 -39 181
rect 39 147 45 181
rect 113 147 119 181
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
rect -119 -181 -113 -147
rect -45 -181 -39 -147
rect 39 -181 45 -147
rect 113 -181 119 -147
<< viali >>
rect -113 147 -103 181
rect -103 147 -55 181
rect -55 147 -45 181
rect 45 147 55 181
rect 55 147 103 181
rect 103 147 113 181
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect -113 -181 -103 -147
rect -103 -181 -55 -147
rect -55 -181 -45 -147
rect 45 -181 55 -147
rect 55 -181 103 -147
rect 103 -181 113 -147
<< metal1 >>
rect -125 181 -33 187
rect -125 147 -113 181
rect -45 147 -33 181
rect -125 141 -33 147
rect 33 181 125 187
rect 33 147 45 181
rect 113 147 125 181
rect 33 141 125 147
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect -125 -147 -33 -141
rect -125 -181 -113 -147
rect -45 -181 -33 -147
rect -125 -187 -33 -181
rect 33 -147 125 -141
rect 33 -181 45 -147
rect 113 -181 125 -147
rect 33 -187 125 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 2 diffcov 100 polycov 70 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
