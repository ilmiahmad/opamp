magic
tech sky130A
magscale 1 2
timestamp 1729232295
<< nmos >>
rect -189 -131 -29 69
rect 29 -131 189 69
<< ndiff >>
rect -247 57 -189 69
rect -247 -119 -235 57
rect -201 -119 -189 57
rect -247 -131 -189 -119
rect -29 57 29 69
rect -29 -119 -17 57
rect 17 -119 29 57
rect -29 -131 29 -119
rect 189 57 247 69
rect 189 -119 201 57
rect 235 -119 247 57
rect 189 -131 247 -119
<< ndiffc >>
rect -235 -119 -201 57
rect -17 -119 17 57
rect 201 -119 235 57
<< poly >>
rect -189 141 -29 157
rect -189 107 -173 141
rect -45 107 -29 141
rect -189 69 -29 107
rect 29 141 189 157
rect 29 107 45 141
rect 173 107 189 141
rect 29 69 189 107
rect -189 -157 -29 -131
rect 29 -157 189 -131
<< polycont >>
rect -173 107 -45 141
rect 45 107 173 141
<< locali >>
rect -189 107 -173 141
rect -45 107 -29 141
rect 29 107 45 141
rect 173 107 189 141
rect -235 57 -201 73
rect -235 -135 -201 -119
rect -17 57 17 73
rect -17 -135 17 -119
rect 201 57 235 73
rect 201 -135 235 -119
<< viali >>
rect -173 107 -45 141
rect 45 107 173 141
rect -235 -119 -201 57
rect -17 -119 17 57
rect 201 -119 235 57
<< metal1 >>
rect -185 141 -33 147
rect -185 107 -173 141
rect -45 107 -33 141
rect -185 101 -33 107
rect 33 141 185 147
rect 33 107 45 141
rect 173 107 185 141
rect 33 101 185 107
rect -241 57 -195 69
rect -241 -119 -235 57
rect -201 -119 -195 57
rect -241 -131 -195 -119
rect -23 57 23 69
rect -23 -119 -17 57
rect 17 -119 23 57
rect -23 -131 23 -119
rect 195 57 241 69
rect 195 -119 201 57
rect 235 -119 241 57
rect 195 -131 241 -119
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
