magic
tech sky130A
magscale 1 2
timestamp 1729261955
<< nwell >>
rect -176 -104 822 2789
<< nsubdiff >>
rect -140 2719 -80 2753
rect 726 2719 786 2753
rect -140 2693 -106 2719
rect 752 2693 786 2719
rect -140 -34 -106 -8
rect 752 -34 786 -8
rect -140 -68 -80 -34
rect 726 -68 786 -34
<< nsubdiffcont >>
rect -80 2719 726 2753
rect -140 -8 -106 2693
rect 752 -8 786 2693
rect -80 -68 726 -34
<< poly >>
rect -56 2681 36 2697
rect -56 2647 -40 2681
rect -6 2647 36 2681
rect -56 2631 36 2647
rect 6 2626 36 2631
rect 610 2681 702 2697
rect 610 2647 652 2681
rect 686 2647 702 2681
rect 610 2632 702 2647
rect 610 2626 640 2632
rect -56 1981 36 1997
rect 94 1996 294 2104
rect -56 1947 -40 1981
rect -6 1947 36 1981
rect -56 1931 36 1947
rect 6 1926 36 1931
rect 610 1981 702 1997
rect 610 1947 652 1981
rect 686 1947 702 1981
rect 610 1932 702 1947
rect 610 1926 640 1932
rect 94 1296 552 1404
rect 6 753 36 782
rect -56 738 36 753
rect -56 704 -40 738
rect -6 704 36 738
rect 610 757 640 775
rect 610 742 702 757
rect 610 708 652 742
rect 686 708 702 742
rect -56 688 36 704
rect 352 596 552 704
rect 610 692 702 708
rect 6 53 36 78
rect -56 38 36 53
rect -56 4 -40 38
rect -6 4 36 38
rect -56 -12 36 4
rect 610 57 640 75
rect 610 42 702 57
rect 610 8 652 42
rect 686 8 702 42
rect 610 -8 702 8
<< polycont >>
rect -40 2647 -6 2681
rect 652 2647 686 2681
rect -40 1947 -6 1981
rect 652 1947 686 1981
rect -40 704 -6 738
rect 652 708 686 742
rect -40 4 -6 38
rect 652 8 686 42
<< locali >>
rect -140 2719 -80 2753
rect 726 2719 786 2753
rect -140 2693 -106 2719
rect 752 2693 786 2719
rect -56 2647 -40 2681
rect -6 2647 10 2681
rect 636 2647 652 2681
rect 686 2647 702 2681
rect -40 2604 -6 2647
rect 652 2604 686 2647
rect -56 1947 -40 1981
rect -6 1947 10 1981
rect 636 1947 652 1981
rect 686 1947 702 1981
rect -40 1904 -6 1947
rect 652 1904 686 1947
rect -40 738 -6 800
rect 652 742 686 796
rect -56 704 -40 738
rect -6 704 10 738
rect 636 708 652 742
rect 686 708 702 742
rect -40 38 -6 102
rect 652 42 686 98
rect -56 4 -40 38
rect -6 4 10 38
rect 636 8 652 42
rect 686 8 702 42
rect -140 -34 -106 -8
rect 752 -34 786 -8
rect -140 -68 -80 -34
rect 726 -68 786 -34
<< viali >>
rect 652 2719 686 2753
rect -40 2647 -6 2681
rect 652 2647 686 2681
rect -40 1947 -6 1981
rect 652 1947 686 1981
rect -40 704 -6 738
rect 652 708 686 742
rect -40 4 -6 38
rect 652 8 686 42
rect -40 -68 -6 -34
<< metal1 >>
rect 640 2753 698 2759
rect 640 2719 652 2753
rect 686 2719 698 2753
rect -52 2681 6 2687
rect -52 2647 -40 2681
rect -6 2647 6 2681
rect -52 2641 6 2647
rect 640 2681 698 2719
rect 640 2647 652 2681
rect 686 2647 698 2681
rect 640 2641 698 2647
rect -46 2600 0 2641
rect 646 2600 692 2641
rect -46 2588 88 2600
rect -59 2212 -49 2588
rect 3 2212 88 2588
rect -46 2200 88 2212
rect 300 2158 346 2600
rect 558 2200 692 2600
rect 558 2158 604 2200
rect 300 2114 382 2158
rect 522 2114 604 2158
rect -52 1981 6 1987
rect -52 1947 -40 1981
rect -6 1947 6 1981
rect -52 1941 6 1947
rect -46 1900 0 1941
rect -46 1888 88 1900
rect -46 1512 38 1888
rect 90 1512 100 1888
rect -46 1500 88 1512
rect 42 1242 124 1286
rect 42 1200 88 1242
rect -46 800 88 1200
rect -46 744 0 800
rect -52 738 6 744
rect -52 704 -40 738
rect -6 704 6 738
rect -52 698 6 704
rect 300 586 346 2114
rect 640 1981 698 1987
rect 640 1947 652 1981
rect 686 1947 698 1981
rect 640 1941 698 1947
rect 646 1900 692 1941
rect 558 1500 692 1900
rect 558 1458 604 1500
rect 522 1414 604 1458
rect 558 1188 692 1200
rect 544 812 554 1188
rect 606 812 692 1188
rect 558 800 692 812
rect 646 748 692 800
rect 640 742 698 748
rect 640 708 652 742
rect 686 708 698 742
rect 640 702 698 708
rect 42 542 124 586
rect 264 542 346 586
rect 42 500 88 542
rect -46 100 88 500
rect 300 100 346 542
rect 558 488 692 500
rect 558 112 642 488
rect 694 112 704 488
rect 558 100 692 112
rect -46 44 0 100
rect 646 48 692 100
rect -52 38 6 44
rect -52 4 -40 38
rect -6 4 6 38
rect -52 -34 6 4
rect 640 42 698 48
rect 640 8 652 42
rect 686 8 698 42
rect 640 2 698 8
rect -52 -68 -40 -34
rect -6 -68 6 -34
rect -52 -74 6 -68
<< via1 >>
rect -49 2212 3 2588
rect 38 1512 90 1888
rect 554 812 606 1188
rect 642 112 694 488
<< metal2 >>
rect -49 2588 3 2598
rect -49 2090 3 2212
rect -49 2081 16 2090
rect -49 2020 -45 2081
rect 629 2020 638 2080
rect 698 2020 707 2080
rect -49 2011 16 2020
rect -49 676 3 2011
rect 38 1888 90 1898
rect 38 1372 90 1512
rect 38 1320 606 1372
rect 554 1188 606 1320
rect 554 802 606 812
rect 642 686 694 2020
rect 628 677 694 686
rect -62 616 -53 676
rect 7 616 16 676
rect 690 615 694 677
rect 628 606 694 615
rect 642 488 694 606
rect 642 102 694 112
<< via2 >>
rect -45 2020 16 2081
rect 638 2020 698 2080
rect -53 616 7 676
rect 628 615 690 677
<< metal3 >>
rect -50 2081 704 2086
rect -50 2020 -45 2081
rect 16 2080 704 2081
rect 16 2020 638 2080
rect 698 2020 704 2080
rect -50 2015 704 2020
rect -59 677 695 682
rect -59 676 628 677
rect -59 616 -53 676
rect 7 616 628 676
rect -59 615 628 616
rect 690 615 695 677
rect -59 610 695 615
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729173951
transform 1 0 625 0 1 300
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729173951
transform 1 0 21 0 1 300
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729173951
transform 1 0 21 0 1 2400
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729173951
transform 1 0 21 0 1 1700
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729173951
transform 1 0 21 0 1 1000
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729173951
transform 1 0 625 0 1 2400
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729173951
transform 1 0 625 0 1 1700
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729173951
transform 1 0 625 0 1 1000
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729173951
transform 1 0 323 0 1 300
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729173951
transform 1 0 323 0 1 1000
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729173951
transform 1 0 323 0 1 1700
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729173951
transform 1 0 323 0 1 2400
box -323 -300 323 300
<< labels >>
flabel metal1 669 2707 669 2707 0 FreeSans 160 0 0 0 vdd
port 1 nsew
flabel metal2 81 1344 81 1344 0 FreeSans 160 0 0 0 d1
port 2 nsew
flabel metal1 581 1442 581 1442 0 FreeSans 160 0 0 0 d2
port 3 nsew
flabel metal2 669 1381 669 1381 0 FreeSans 160 0 0 0 d5
port 4 nsew
flabel metal2 68 1380 68 1380 0 FreeSans 160 0 0 0 d1
flabel metal1 584 1468 584 1468 0 FreeSans 160 0 0 0 d2
flabel metal2 668 1336 668 1336 0 FreeSans 160 0 0 0 d5
flabel metal1 672 2610 672 2610 0 FreeSans 160 0 0 0 vdd
<< end >>
