magic
tech sky130A
magscale 1 2
timestamp 1729197478
<< nwell >>
rect -223 -200 223 200
<< pmos >>
rect -129 -100 -29 100
rect 29 -100 129 100
<< pdiff >>
rect -187 88 -129 100
rect -187 -88 -175 88
rect -141 -88 -129 88
rect -187 -100 -129 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 129 88 187 100
rect 129 -88 141 88
rect 175 -88 187 88
rect 129 -100 187 -88
<< pdiffc >>
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
<< poly >>
rect -112 181 -46 197
rect -112 164 -96 181
rect -129 147 -96 164
rect -62 164 -46 181
rect 46 181 112 197
rect 46 164 62 181
rect -62 147 -29 164
rect -129 100 -29 147
rect 29 147 62 164
rect 96 164 112 181
rect 96 147 129 164
rect 29 100 129 147
rect -129 -147 -29 -100
rect -129 -164 -96 -147
rect -112 -181 -96 -164
rect -62 -164 -29 -147
rect 29 -147 129 -100
rect 29 -164 62 -147
rect -62 -181 -46 -164
rect -112 -197 -46 -181
rect 46 -181 62 -164
rect 96 -164 129 -147
rect 96 -181 112 -164
rect 46 -197 112 -181
<< polycont >>
rect -96 147 -62 181
rect 62 147 96 181
rect -96 -181 -62 -147
rect 62 -181 96 -147
<< locali >>
rect -175 88 -141 104
rect -175 -104 -141 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 141 88 175 104
rect 141 -104 175 -88
<< viali >>
rect -113 147 -96 181
rect -96 147 -62 181
rect -62 147 -45 181
rect 45 147 62 181
rect 62 147 96 181
rect 96 147 113 181
rect -175 -88 -141 88
rect -17 -88 17 88
rect 141 -88 175 88
rect -113 -181 -96 -147
rect -96 -181 -62 -147
rect -62 -181 -45 -147
rect 45 -181 62 -147
rect 62 -181 96 -147
rect 96 -181 113 -147
<< metal1 >>
rect -125 181 -33 187
rect -125 147 -113 181
rect -45 147 -33 181
rect -125 141 -33 147
rect 33 181 125 187
rect 33 147 45 181
rect 113 147 125 181
rect 33 141 125 147
rect -181 88 -135 100
rect -181 -88 -175 88
rect -141 -88 -135 88
rect -181 -100 -135 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 135 88 181 100
rect 135 -88 141 88
rect 175 -88 181 88
rect 135 -100 181 -88
rect -125 -147 -33 -141
rect -125 -181 -113 -147
rect -45 -181 -33 -147
rect -125 -187 -33 -181
rect 33 -147 125 -141
rect 33 -181 45 -147
rect 113 -181 125 -147
rect 33 -187 125 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 2 diffcov 100 polycov 20 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
