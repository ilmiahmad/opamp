magic
tech sky130A
magscale 1 2
timestamp 1729262064
<< psubdiff >>
rect -190 207 -130 241
rect 1018 207 1078 241
rect -190 181 -156 207
rect 1044 181 1078 207
rect -190 -1208 -156 -1186
rect 1044 -1208 1078 -1186
rect -190 -1242 -130 -1208
rect 1018 -1242 1078 -1208
<< psubdiffcont >>
rect -130 207 1018 241
rect -190 -1186 -156 181
rect 1044 -1186 1078 181
rect -130 -1242 1018 -1208
<< poly >>
rect -106 -338 -40 -334
rect -106 -350 -14 -338
rect -106 -384 -90 -350
rect -56 -384 -14 -350
rect -106 -400 -14 -384
rect 902 -350 994 -334
rect 902 -384 944 -350
rect 978 -384 994 -350
rect 902 -400 994 -384
rect 158 -600 730 -400
rect -106 -616 -14 -600
rect -106 -650 -90 -616
rect -56 -650 -14 -616
rect -106 -666 -14 -650
rect 902 -616 994 -600
rect 902 -650 944 -616
rect 978 -650 994 -616
rect 902 -666 994 -650
<< polycont >>
rect -90 -384 -56 -350
rect 944 -384 978 -350
rect -90 -650 -56 -616
rect 944 -650 978 -616
<< locali >>
rect -190 207 -130 241
rect 1018 207 1078 241
rect -190 181 -156 207
rect 1044 181 1078 207
rect -90 -350 -56 -316
rect 944 -350 978 -316
rect -106 -384 -90 -350
rect -56 -384 -40 -350
rect 928 -384 944 -350
rect 978 -384 994 -350
rect -106 -650 -90 -616
rect -56 -650 -40 -616
rect 928 -650 944 -616
rect 978 -650 994 -616
rect -90 -684 -56 -650
rect 944 -684 978 -650
rect -190 -1208 -156 -1186
rect 1044 -1208 1078 -1186
rect -190 -1242 -130 -1208
rect 1018 -1242 1078 -1208
<< viali >>
rect 364 207 410 241
rect -90 -300 -56 76
rect -2 -300 32 76
rect 112 -300 146 76
rect 370 -300 404 76
rect 484 -300 518 76
rect 742 -300 776 76
rect 856 -300 890 76
rect 944 -300 978 76
rect -90 -384 -56 -350
rect 174 -384 342 -350
rect 944 -384 978 -350
rect -90 -650 -56 -616
rect 546 -650 714 -616
rect 944 -650 978 -616
rect -90 -1076 -56 -700
rect -2 -1076 32 -700
rect 112 -1076 146 -700
rect 370 -1076 404 -700
rect 484 -1076 518 -700
rect 742 -1076 776 -700
rect 856 -1076 890 -700
rect 944 -1076 978 -700
rect 478 -1242 524 -1208
<< metal1 >>
rect 351 197 361 249
rect 413 197 423 249
rect -96 76 152 88
rect 364 76 410 88
rect 478 76 524 88
rect 736 76 984 88
rect -96 -300 -90 76
rect -56 -300 -2 76
rect 32 -300 112 76
rect 146 -300 152 76
rect 351 -300 361 76
rect 413 -300 423 76
rect 465 -300 475 76
rect 527 -300 537 76
rect 736 -300 742 76
rect 776 -300 856 76
rect 890 -300 944 76
rect 978 -300 984 76
rect -96 -312 152 -300
rect 364 -312 410 -300
rect 478 -312 524 -300
rect 736 -312 984 -300
rect -96 -344 -50 -312
rect 106 -344 152 -312
rect -102 -350 -44 -344
rect -102 -384 -90 -350
rect -56 -384 -44 -350
rect -102 -390 -44 -384
rect 106 -350 354 -344
rect 106 -384 174 -350
rect 342 -384 354 -350
rect 106 -390 354 -384
rect 788 -472 844 -312
rect 938 -344 984 -312
rect 932 -350 990 -344
rect 932 -384 944 -350
rect 978 -384 990 -350
rect 932 -390 990 -384
rect 44 -528 844 -472
rect -102 -616 -44 -610
rect -102 -650 -90 -616
rect -56 -650 -44 -616
rect -102 -656 -44 -650
rect -96 -688 -50 -656
rect 44 -688 100 -528
rect 534 -616 782 -610
rect 534 -650 546 -616
rect 714 -650 782 -616
rect 534 -656 782 -650
rect 932 -616 990 -610
rect 932 -650 944 -616
rect 978 -650 990 -616
rect 932 -656 990 -650
rect 736 -688 782 -656
rect 944 -688 978 -656
rect -96 -700 152 -688
rect 364 -700 410 -688
rect 478 -700 524 -688
rect 736 -700 984 -688
rect -96 -1076 -90 -700
rect -56 -1076 -2 -700
rect 32 -1076 112 -700
rect 146 -1076 152 -700
rect 351 -1076 361 -700
rect 413 -1076 423 -700
rect 465 -1076 475 -700
rect 527 -1076 537 -700
rect 736 -1076 742 -700
rect 776 -1076 856 -700
rect 890 -1076 944 -700
rect 978 -1076 984 -700
rect -96 -1088 152 -1076
rect 364 -1088 410 -1076
rect 478 -1089 524 -1076
rect 736 -1088 984 -1076
rect 465 -1250 475 -1198
rect 527 -1250 537 -1198
<< via1 >>
rect 361 241 413 249
rect 361 207 364 241
rect 364 207 410 241
rect 410 207 413 241
rect 361 197 413 207
rect 361 -300 370 76
rect 370 -300 404 76
rect 404 -300 413 76
rect 475 -300 484 76
rect 484 -300 518 76
rect 518 -300 527 76
rect 361 -1076 370 -700
rect 370 -1076 404 -700
rect 404 -1076 413 -700
rect 475 -1076 484 -700
rect 484 -1076 518 -700
rect 518 -1076 527 -700
rect 475 -1208 527 -1198
rect 475 -1242 478 -1208
rect 478 -1242 524 -1208
rect 524 -1242 527 -1208
rect 475 -1250 527 -1242
<< metal2 >>
rect 361 249 413 259
rect 361 76 413 197
rect 361 -474 413 -300
rect 473 76 529 86
rect 473 -310 529 -300
rect 361 -526 527 -474
rect 359 -700 415 -690
rect 359 -1086 415 -1076
rect 475 -700 527 -526
rect 475 -1198 527 -1076
rect 475 -1260 527 -1250
<< via2 >>
rect 473 -300 475 76
rect 475 -300 527 76
rect 527 -300 529 76
rect 359 -1076 361 -700
rect 361 -1076 413 -700
rect 413 -1076 415 -700
<< metal3 >>
rect 463 76 539 81
rect 463 -300 473 76
rect 529 -300 539 76
rect 463 -461 539 -300
rect 349 -537 539 -461
rect 349 -700 425 -537
rect 349 -1076 359 -700
rect 415 -1076 425 -700
rect 349 -1081 425 -1076
use sky130_fd_pr__nfet_01v8_Q6XT6P  sky130_fd_pr__nfet_01v8_Q6XT6P_0
timestamp 1729185943
transform 1 0 444 0 1 -112
box -344 -288 344 288
use sky130_fd_pr__nfet_01v8_Q6XT6P  sky130_fd_pr__nfet_01v8_Q6XT6P_1
timestamp 1729185943
transform 1 0 444 0 1 -888
box -344 -288 344 288
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_0
timestamp 1729184572
transform 1 0 -29 0 1 -888
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_1
timestamp 1729184572
transform 1 0 917 0 1 -888
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_2
timestamp 1729184572
transform 1 0 -29 0 1 -112
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_TC9PLT  sky130_fd_pr__nfet_01v8_TC9PLT_4
timestamp 1729184572
transform 1 0 917 0 1 -112
box -73 -226 73 226
<< labels >>
flabel space 258 -107 258 -107 0 FreeSans 160 0 0 0 m3
flabel space 246 -937 246 -937 0 FreeSans 160 0 0 0 m4
flabel viali 503 -1003 503 -1003 0 FreeSans 160 0 0 0 m3
flabel viali 511 -119 511 -119 0 FreeSans 160 0 0 0 m4
flabel metal2 383 141 383 141 0 FreeSans 160 0 0 0 vgnd
port 1 nsew
flabel metal3 388 -647 388 -647 0 FreeSans 160 0 0 0 rs
port 2 nsew
flabel metal1 127 -368 127 -368 0 FreeSans 160 0 0 0 d3
port 3 nsew
flabel metal1 813 -500 813 -500 0 FreeSans 160 0 0 0 d4
port 4 nsew
flabel metal1 814 -420 814 -420 0 FreeSans 160 0 0 0 d4
flabel metal1 126 -338 126 -338 0 FreeSans 160 0 0 0 d3
flabel metal3 384 -624 384 -624 0 FreeSans 160 0 0 0 rs
flabel metal2 386 172 386 172 0 FreeSans 160 0 0 0 vgnd
<< end >>
